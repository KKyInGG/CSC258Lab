
module combine(SW,KEY,state);
	input [9:0] SW;
	input [3:0] KEY;
	output [7:0] fx;
	output [6:0] fy;
	output [2:0] fc;
	
	wire x1,y1,c1,start1;
	controller c1(
		.rset(KEY[0]),
		.clk(KEY[2]),
		.go(KEY[3]),
		.draw(KEY[1]),
		.lx(x1),
		.ly(y1),
		.lc(c1),
		.start(start1),
	);
	
	datapath d1(
		.colour(SW[7:9]), 
		.clk(KEY[2]), 
		.loc_in(SW[6:0]), 
		.en_x(x1), 
		.en_y(y1), 
		.en_c(c1), 
		.en_ix(start1), 
		.r_set(KEY[0]), 
		.sx(fx), 
		.sy(fy), 
		.sc(fc)
		);

module controller (rset, clk, go, draw, lx, ly, lc, start, state );
	input rset,clk,go,draw;
	output reg lx,ly,lc,start;
	output [2:0] state;
	
	reg [2:0] current,next;
	
	localparam Load_x_wait = 3'd0,
				  Load_x = 3'd1,
				  Load_y_wait = 3'd2,
				  Load_y = 3'd3,
				  Draw = 3'd4;
	
	 always @(*)
		begin
			case(current)
				Load_x_wait: next = go ? Load_x : Load_x_wait;
				Load_x : next = go ? Load_x : Load_y_wait;
				Load_y_wait : next = go ? Load_y_wait : Load_y;
				Load_y : next = draw ? Load_y : Draw;
				Draw : next = Load_x_wait;
				default: next = Load_x_wait;
			endcase
		end
		
	
	  always @(*) 
		begin
			lx = 1'b0;
			ly = 1'b0;
			lc = 1'b0;
			start = 1'b0;
			
			case(current)
				Load_x_wait: lx = 1'b1;
				Load_y_wait:
					begin
						ly = 1'b1;
						lc = 1'b1;
					end
				Draw: start = 1'b1;
			endcase
	  end
	  
	  always @(posedge clk)
			begin
				if(!rset)
					current <= Load_x_wait;
				else
					current <= next;
			end
		assign state = current;
endmodule

				
	
module datapath (colour, clk, loc_in, en_x, en_y, en_c, en_ix, r_set, sx, sy, sc );
		input [6:0] loc_in;
		input [2:0] colour;
		input clk,r_set;
		input en_x, en_y, en_c, en_ix;
		reg en_iy;
		output [7:0] sx;
		output [6:0]sy;
		output [2:0] sc;
		
		reg [7:0] x;
		reg [6:0] y;
		reg [2:0] c;	
		
		always @(posedge clk)
			begin
				if(!r_set)
					begin
						x <= 8'd0;
						y <= 7'd0;
						c <= 3'd0;
					end
				else
					begin
						if(en_x)
							x <= {1'b0, loc_in};
						if(en_y)
							y <= {loc_in};
						if (en_c)
							c <= colour;
					end
			end
	  
	  reg [1:0] ix;
	  reg [1:0] iy;
			
	  always @(posedge clk)
			begin
				if(!r_set)
					begin
						ix <= 2'd0;
						iy <= 2'd0;
					end
				if(en_ix)
					if (ix == 2'b11)
					   begin
							ix <= 2'b00;
							en_iy <= 1'b1;
						end
					else
						begin
							ix <= ix + 2'b01;
							en_iy <= 1'b0;
						end
			end
			
		  always @(posedge clk)
			begin
				if(!r_set)
					begin
						ix <= 2'd0;
						iy <= 2'd0;
					end
				if(en_iy)
					if (iy == 2'b11)
					   begin
							iy <= 2'b00;
						end
					else
						iy <= iy + 2'b01;
			end
			
			assign sx = x + ix;
			assign sy = y + iy;
			assign sc = c;
			
endmodule
